module ALU (
	input[15:0] data1,
	input[15:0] data2,
	output[15:0] zero, // TODO check if this is 16 bit
	output[15:0] result,
	input[2:0] ALU_control_output
);
	//TODO
endmodule