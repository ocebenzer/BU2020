module Adder()