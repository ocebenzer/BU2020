module RegisterMux()