`timescale 1ns/1ns

module Memory(
	input clk,
	input[11:0] address_bus,
	output[15:0] data_bus,
	input[15:0] incoming_data_bus,
	input write_mode,
	input[11:0] Instruction_addressbus,
	output[15:0] Instruction_databus,
	input doubleRead,
	input doubleWrite
	);

	// 4KB Memory, 4x1KB modules, first module is instruction module, rest 3 are data modules
	reg[511:0][15:0] data_instruction = 8192'hD000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000D000;
	reg[511:0][15:0] data1 = 8192'h10001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000;
	reg[511:0][15:0] data2 = 8192'h20002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000200020002000;
	reg[511:0][15:0] data3 = 8192'h30003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000300030003000;
	
	initial begin
	//Instruction Initialization

 		//jump to decimal 400 instructions, pass the next 15 instructions
		data_instruction[0] = 16'hF190;
/*
		//0000 010 011 100 XXX, 04E0h Add R010 R011 R100
		data_instruction[5] = 16'h04E0;
		//0001 010 011 000110, 14C6h Add R010 R011 memory(BA+"6")
		data_instruction[10] = 16'h14C6;
		//0010 010 011 100 XXX, 24E0h Sub R010 R011 R100
		data_instruction[20] = 16'h24E0;
		//0011 010 011 000110, 34C6h Addi R010 R011  "6"
		data_instruction[30] = 16'h34C6;
		//0100 010 011 100 XXX, 44E0h Mul R010 R011 R100
		data_instruction[40] = 16'h44E0;
		//0101 010 011 100 XXX, 54E0h And R010 R011 R100
		data_instruction[50] = 16'h54E0;
		//0110 010 000001001, 6409h Sll R010 "9"
		data_instruction[60] = 16'h6409;
		//0111 010 000001001, 7409h Lw R010 "9"
		data_instruction[70] = 16'h7409;
		//1000 010 000001001, 8409h Lwi R010 "9"
		data_instruction[80] = 16'h8409;
		//1001 010 000001001, 9409h Sw R010 "9"
		data_instruction[90] = 16'h9409;
		//1010 010 000001001, A409h Swi R010 "9"
		data_instruction[100] = 16'hA409;
		//1011 010 XXXXXXXXX, B400h CLR R010
		data_instruction[110] = 16'hB400;
		//1100 010 000001001, C409h Mov R010 "9"
		data_instruction[120] = 16'hC409;
		//1101 XXX 011 100 XXX, D0E0h CMP R011 R100
		data_instruction[130] = 16'hD0E0;
		//1110 000100000000, E00Ch Bne "Pc + 2x256"
		data_instruction[140] = 16'hE100;
		//1111 000000000000, F4ECh Jmp "2x0"
		data_instruction[150] = 16'hF000;
*/
	// decimal 400 instructions start here

		//0000 011 010 001 XXX, 04E0h Add 011 010 001
		data_instruction[200] = 16'h0688;
		//0010 100 010 011 XXX, 24E0h Sub R100 R011 R010
		data_instruction[210] = 16'h2898;
		//0011 101 100 100000, 34C6h Addi R101 R100  "32"
		data_instruction[220] = 16'h3B20;
		//0100 110 110 000 XXX, 44E0h Mul R110 R110 R000
		data_instruction[230] = 16'h4D80;
		//0101 111 100 110 XXX, 54E0h And R111 R100 R110
		data_instruction[240] = 16'h5F30;
		//0110 111 000000001, 6409h Sll R111 "1"
		data_instruction[250] = 16'h6E01;
		//0111 010 000001001, 7409h Lw R010 "BA+2x9"
		data_instruction[260] = 16'h7409;
		//1001 010 000001010, 9409h Sw R010 "BA+2x10"
		data_instruction[270] = 16'h940A;
		//1011 010 XXXXXXXXX, B400h CLR R010
		data_instruction[280] = 16'hB400;
		//1100 010 000001001, C409h Mov R010 "9"
		data_instruction[290] = 16'hC409;

		
		//1000 111 000110000, 8409h Lwi R111 "48"
		data_instruction[350] = 16'h8E30;
		//0011 111 111 000001, 34C6h Addi R111 R111  "1"
		data_instruction[355] = 16'h3FC1;
		//1010 111 000110001, A409h Swi R111 "49"
		data_instruction[360] = 16'hAE31;

		/*
		data_instruction[200] = 16'hD050; // CMP R010 R001
		data_instruction[201] = 16'hEFFF; // Bne (Pc + 2 x "-1")
		*/

	//The ultimate script

		data_instruction[400] = 16'hCEFF;	// Mov $111 0xFF
		data_instruction[405] = 16'h6E04;	// Sll $111 "4"
		data_instruction[410] = 16'h31C0;	// Addi $000 $111 0x0 - 0011 001 111 001010
		data_instruction[411] = 16'h33CE;	// Addi $001 $111 0xE - 0011 000 111 001111
		data_instruction[412] = 16'h35C0;	// Addi $010 $111 0x0 - 0011 010 111 000000
		data_instruction[415] = 16'h3002;	// Addi $000 $000 "2" - 0011 000 000 000001 *LOOP
		data_instruction[420] = 16'h9400;	// Sw $010 "0"
		data_instruction[425] = 16'hD008;	// Cmp $000 $001 - D xxx 000 001 xxx
		data_instruction[426] = 16'hEFF5;	// Bne 2 x "-11" - 1110 0x-11
		
	// Memory Initialization
		data1[9] <= 16'h0018;
		data1[48] <= 16'h07FE;
		data1[49] <= 16'h07FF;
		data1[510] <= 16'hcccc;
		data1[511] <= 16'hbbbb;

		/*
		12 bit adres
		2 bit -> blok
		9 bit -> data
		1 bit -> dont care
		*/
	end

	// Read Data
	reg[15:0] data_bus_init_read, data_bus_final_read;
	assign data_bus = data_bus_final_read;
	always @ * begin
		// Initial read
		case(address_bus[11:10])
			2'b00: data_bus_init_read <= data_instruction[address_bus[9:1]];
			2'b01: data_bus_init_read <= data1[address_bus[9:1]];
			2'b10: data_bus_init_read <= data2[address_bus[9:1]];
			2'b11: data_bus_init_read <= data3[address_bus[9:1]];
		endcase

		case (doubleRead)
			1'b1: begin
				case(data_bus_init_read[11:10])
					2'b00: data_bus_final_read <= data_instruction[data_bus_init_read[9:1]];
					2'b01: data_bus_final_read <= data1[data_bus_init_read[9:1]];
					2'b10: data_bus_final_read <= data2[data_bus_init_read[9:1]];
					2'b11: data_bus_final_read <= data3[data_bus_init_read[9:1]];
				endcase
			end
			default: data_bus_final_read <= data_bus_init_read;
		endcase
	end

	// Write Data
	always@(posedge clk) begin
		case (write_mode)
			1'b1: begin
				case (doubleWrite)
					1'b1: begin
						case(data_bus_init_read[11:10])
							2'b00: data_instruction[data_bus_init_read[9:1]] <= incoming_data_bus;
							2'b01: data1[data_bus_init_read[9:1]] <= incoming_data_bus;
							2'b10: data2[data_bus_init_read[9:1]] <= incoming_data_bus;
							2'b11: data3[data_bus_init_read[9:1]] <= incoming_data_bus;
						endcase
					end
					default: begin
						case(address_bus[11:10])
							2'b00: data_instruction[address_bus[9:1]] <= incoming_data_bus;
							2'b01: data1[address_bus[9:1]] <= incoming_data_bus;
							2'b10: data2[address_bus[9:1]] <= incoming_data_bus;
							2'b11: data3[address_bus[9:1]] <= incoming_data_bus;
						endcase
					end
				endcase
			end
		endcase
	end

	// Read Instruction
	assign Instruction_databus =
		(Instruction_addressbus[11:10] == 2'b00) ? data_instruction[Instruction_addressbus[9:1]]
		: (Instruction_addressbus[11:10] == 2'b01) ? data1[Instruction_addressbus[9:1]]
		: (Instruction_addressbus[11:10] == 2'b10) ? data2[Instruction_addressbus[9:1]]
													: data3[Instruction_addressbus[9:1]];
endmodule